LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY leddec IS
	PORT (
		data : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		anode : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		seg : OUT STD_LOGIC_VECTOR (0 TO 6)
	);
END leddec;

ARCHITECTURE Behavioral OF leddec IS
BEGIN
	-- Turn on segments corresponding to 4-bit data word
	seg <= "0000001" WHEN data = "1111" ELSE --0
	       "1001111" WHEN data = "1110" ELSE --1
	       "0010010" WHEN data = "1101" ELSE --2
	       "0000110" WHEN data = "1100" ELSE --3
	       "1001100" WHEN data = "1011" ELSE --4
	       "0100100" WHEN data = "1010" ELSE --5
	       "0100000" WHEN data = "1001" ELSE --6
	       "0001111" WHEN data = "1000" ELSE --7
	       "0000000" WHEN data = "0111" ELSE --8
	       "0000100" WHEN data = "0110" ELSE --9
	       "0001000" WHEN data = "0101" ELSE --A
	       "1100000" WHEN data = "0100" ELSE --B
	       "0110001" WHEN data = "0011" ELSE --C
	       "1000010" WHEN data = "0010" ELSE --D
	       "0110000" WHEN data = "0001" ELSE --E
	       "0111000" WHEN data = "0000" ELSE --F
	       "1111111";
	-- Turn on anode of 7-segment display addressed by 2-bit digit selector dig
	anode <= "1111";
END Behavioral;
